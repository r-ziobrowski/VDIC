class shape;
	real width_1;
	real width_2;
	real height;
	
	function new();
	endfunction
	
	function real get_area();
	endfunction
	
	function void print();
	endfunction
	
endclass
